`include "uvm_macros.svh"
import uvm_pkg::*;

package Leds_7_test_pkg;
    
    `include "../testbench/uart_sequence_item.svh"
    `include "../testbench/uart_agent.svh"

    `include "../testbench/base_test.svh"
    
endpackage