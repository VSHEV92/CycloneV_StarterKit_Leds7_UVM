// интерфейс сброса блока
  	interface reset_intf();

	    logic resetn = 0;
	    
	 endinterface : reset_intf